// https://www.youtube.com/watch?v=Q-UeYEpwXXU

// Output: [0, 180]

module angles (
    input  logic [1:0] x,
    input  logic [1:0] y,
    output logic [7:0] tan,
    output logic [7:0] cos
);

    real 
endmodule
